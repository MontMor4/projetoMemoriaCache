library verilog;
use verilog.vl_types.all;
entity teste_memoriaCache is
end teste_memoriaCache;
